/*------------------------------------------------------------------------------
 * File          : mmg_driver.sv
 * Project       : RTL
 * Author        : eposmk
 * Creation date : May 17, 2025
 * Description   :
 *------------------------------------------------------------------------------*/

class mmg_driver extends uvm_driver#(mmg_trans);
	`uvm_component_utils(mmg_driver)

	virtual mmg_if vif;
	
	uvm_analysis_port#(mmg_trans) ap;

	// Constructor
	function new(string name = "mmg_driver", uvm_component parent = null);
	  super.new(name, parent);
	  ap = new("ap", this);
	endfunction

	// Grab virtual interface
	virtual function void build_phase(uvm_phase phase);
	  super.build_phase(phase);
	  if (!uvm_config_db#(virtual mmg_if)::get(this, "", "vif", vif)) begin
		`uvm_fatal(get_type_name(), "Virtual interface not found")
	  end
	endfunction

	// Main driver loop
	virtual task run_phase(uvm_phase phase);
		mmg_trans tr;

	  wait (!vif.rst);
	  @(posedge vif.clk);
	  
	  forever begin
		  #1ns
		seq_item_port.get_next_item(tr);
		
		vif.enable <= tr.enable;
		vif.pixel  <= tr.pixel;
		vif.last_in_frame   <= tr.last_in_frame;
		vif.wr_background <= tr.wr_background;
		vif.threshold <= tr.threshold;
		ap.write(tr);
		@(posedge vif.clk);

		seq_item_port.item_done();
	  end

	endtask

  endclass
